module NextStateGenerator( // @[:@3.2]
  input   clock, // @[:@4.4]
  input   reset, // @[:@5.4]
  input   io_input_0, // @[:@6.4]
  input   io_input_1, // @[:@6.4]
  input   io_input_2, // @[:@6.4]
  input   io_input_3, // @[:@6.4]
  input   io_input_4, // @[:@6.4]
  input   io_input_5, // @[:@6.4]
  input   io_input_6, // @[:@6.4]
  input   io_input_7, // @[:@6.4]
  input   io_presentState, // @[:@6.4]
  output  io_nextState // @[:@6.4]
);
  wire [1:0] _T_35; // @[NextStateGenerator.scala 10:58:@8.4]
  wire [1:0] _T_36; // @[NextStateGenerator.scala 10:58:@9.4]
  wire [2:0] _T_37; // @[NextStateGenerator.scala 10:58:@10.4]
  wire [1:0] _T_38; // @[NextStateGenerator.scala 10:58:@11.4]
  wire [1:0] _T_39; // @[NextStateGenerator.scala 10:58:@12.4]
  wire [2:0] _T_40; // @[NextStateGenerator.scala 10:58:@13.4]
  wire [3:0] _T_41; // @[NextStateGenerator.scala 10:58:@14.4]
  wire  _T_43; // @[NextStateGenerator.scala 13:33:@15.4]
  wire  _T_45; // @[NextStateGenerator.scala 13:79:@16.4]
  assign _T_35 = io_input_0 + io_input_1; // @[NextStateGenerator.scala 10:58:@8.4]
  assign _T_36 = io_input_2 + io_input_3; // @[NextStateGenerator.scala 10:58:@9.4]
  assign _T_37 = _T_35 + _T_36; // @[NextStateGenerator.scala 10:58:@10.4]
  assign _T_38 = io_input_4 + io_input_5; // @[NextStateGenerator.scala 10:58:@11.4]
  assign _T_39 = io_input_6 + io_input_7; // @[NextStateGenerator.scala 10:58:@12.4]
  assign _T_40 = _T_38 + _T_39; // @[NextStateGenerator.scala 10:58:@13.4]
  assign _T_41 = _T_37 + _T_40; // @[NextStateGenerator.scala 10:58:@14.4]
  assign _T_43 = _T_41 == 4'h2; // @[NextStateGenerator.scala 13:33:@15.4]
  assign _T_45 = _T_41 == 4'h3; // @[NextStateGenerator.scala 13:79:@16.4]
  assign io_nextState = _T_43 ? io_presentState : _T_45; // @[NextStateGenerator.scala 16:16:@18.4]
endmodule
